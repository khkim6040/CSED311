module ALU (
    input [1:0] alu_op,
    input [31:0] alu_in_1,
    input [31:0] alu_in_2,
    output reg [31:0] alu_result,
    output reg alu_bcond
);

    // TODO: Implement ALU operations


endmodule