module ControlUnit (
    input [6:0] part_of_inst,
    output is_jal,
    output is_jalr,
    output branch,
    output mem_read,
    output mem_to_reg,
    output mem_write,
    output alu_src,
    output write_enable,
    output pc_to_reg,
    output is_ecall
);
    // TODO: Microcode for Control Unit

    // TODO: Assign Control signals

    // TODO: Calculate next state

    // TODO: Update state synchronously

    
endmodule