module ALUControlUnit (
    input funct7,
    input[3:0] funct3,
    input[2:0] ALUOp,
    output reg [3:0] alu_op
);

    // TODO: Generate ALU control signal
    

endmodule